///initial memory map
module map_array (input Clk, Reset,

input logic [0:299][4:0] map_in,
output logic [0:299][4:0] map_out 
);



always_ff @(posedge Clk)
// or posedge Reset)
begin
if (Reset)
begin
map_out <= {
 5'h7,	 5'h7,	 5'h7,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,   5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,
 5'h1,	 5'hD,    5'h0,	 5'h2,    5'h0,    5'h0,    5'h2,	 5'h2,	 5'h0,	 5'h2,   5'h0,	 5'h2,	 5'h2,	 5'h0,	 5'h0,	 5'h2,	 5'h2,	 5'h0,	 5'h2,	 5'h1,
 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h2,   5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,
 5'h1,	 5'h2,	 5'h2,	 5'h0,	 5'h0,	 5'h0,	 5'h2,	 5'h2,	 5'h0,	 5'h2,   5'h2,	 5'h2,	 5'h0,	 5'h0,	 5'h2,	 5'h2,	 5'h2,	 5'h0,	 5'h2,	 5'h1,
 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,   5'h2,	 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h0,	 5'h1,
 5'h1,	 5'h0,	 5'h2,	 5'h0,	 5'h0,	 5'h2,	 5'h2,	 5'h2,	 5'h0,	 5'h0,   5'h2,	 5'h2,	 5'h0,	 5'h0,	 5'h2,	 5'h2,	 5'h0,	 5'h0,	 5'h2,	 5'h1,
 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,   5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,
 5'h1,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h2,	 5'h0,	 5'h2,	 5'h0,	 5'h0,   5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h2,	 5'h0,	 5'h0,	 5'h1,
 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h2,   5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h0,	 5'h1,
 5'h1,	 5'h0,	 5'h0,    5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,   5'h2,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h2,	 5'h1,
 5'h1,	 5'h2,	 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,   5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,	 5'h2,	 5'h1,
 5'h1,	 5'h2,	 5'h2,	 5'h2,	 5'h0,	 5'h2,	 5'h2,	 5'h2,	 5'h0,	 5'h2,   5'h2,	 5'h2,	 5'h0,	 5'h0,	 5'h0,	 5'h2,	 5'h0,	 5'h0,	 5'h2,	 5'h1,
 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h2,	 5'h1,	 5'h2,   5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h0,	 5'h1,	 5'h0,    5'h1,
 5'h1,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h0,	 5'h2,	 5'h0,	 5'h0,   5'h2,	 5'h0,	 5'h2,	 5'h0,	 5'h2,	 5'h0,	 5'h2,	 5'h0,	 5'h15,   5'h1,
 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,   5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h1,	 5'h7,	 5'h7,	 5'h7
};
end

else
map_out <=map_in;

end
endmodule 