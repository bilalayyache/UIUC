//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module lab8( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1,
				 output logic [3:0]	LED,
             // VGA Interface 
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK      //SDRAM Clock
                    );
    
    logic Reset_h, Clk;
    logic [7:0] keycode;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            .from_sw_reset(hpi_reset),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),
                            .OTG_RST_N(OTG_RST_N)
    );
     
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     nios_system nios_system(
                             .clk_clk(Clk),         
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w),
                             .otg_hpi_reset_export(hpi_reset)
    );
    
    // Use PLL to generate the 25MHZ VGA_CLK.
    // You will have to generate it on your own in simulation.
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
    
	 // logic for keycode
	 // logic space_on, a_on, s_on, d_on;
	 // keycode_reader keycode_reader_instance(.*);
	 
	 // coordinate for drawing
	 logic[12:0] X, Y;
	 logic		isMario;
	 logic[23:0] ground_dout, stand_dout, cloud_dout, background_dout, L_mountain_dout, S_mountain_dout, tube_1_dout, tube_2_dout, tube_3_dout, castle_dout;
	 
    // TODO: Fill in the connections for the rest of the modules 
    VGA_controller vga_controller_instance(.Clk,
														 .Reset(Reset_h),      
														 .VGA_HS,
														 .VGA_VS,
														 .VGA_CLK,
														 .VGA_BLANK_N,
														 .VGA_SYNC_N,
														 .DrawX(X),
														 .DrawY(Y)       
														);
    
	 logic [12:0] Mario_X_Pos, Mario_Y_Pos, process, Cloud_X_Pos, Cloud_Y_Pos, L_mountain_X_Pos, L_mountain_Y_Pos, S_mountain_X_Pos, S_mountain_Y_Pos;
	 logic [12:0] tube_1_X_Pos, tube_1_Y_Pos, tube_2_X_Pos, tube_2_Y_Pos,tube_3_X_Pos, tube_3_Y_Pos, castle_X_Pos, castle_Y_Pos;
    // Which signal should be frame_clk?
    Mario mario_instance(.Clk,
	                    .Reset(Reset_h),
	                    .frame_clk(VGA_VS),
	                    .DrawX(X), .DrawY(Y),
	                    .is_Mario(isMario),
							  .keycode,
							  .Mario_X_Pos,
							  .Mario_Y_Pos,
							  .process
							 );
    
    color_mapper color_instance(.is_Mario(isMario),
	                             .DrawX(X), .DrawY(Y),
	                             .VGA_R, .VGA_G, .VGA_B,
										  .ground_dout, .stand_dout,
										  .process
										 );
    
	 
	  // we put our background here
	  GROUND ground_instance(.Clk, .read_address((X+process)%32 + 32*(Y%64)), .data_Out(ground_dout));
	  
	  CLOUD cloud_instance(.Clk, .read_address((X-Cloud_X_Pos+process)%64 + 64*((Y-Cloud_Y_Pos)%48)), .data_Out(cloud_dout));
	  
	  LARGE_MOUNTAIN large_mountain_instance(.Clk, .read_address((X-L_mountain_X_Pos+process)%160 + 160*((Y-L_mountain_Y_Pos)%72)), .data_Out(L_mountain_dout));
	
	  MOUNTAIN mountain_instance(.Clk, .read_address((X-S_mountain_X_Pos+process)%64 + 64*((Y-S_mountain_Y_Pos)%32)), .data_Out(S_mountain_dout));
	  
	  TUBE_1 tube_1_instance(.Clk, .read_address((X-tube_1_X_Pos+process)%64 + 64*((Y-tube_1_Y_Pos)%64)), .data_Out(tube_1_dout));
	  TUBE_2 tube_2_instance(.Clk, .read_address((X-tube_2_X_Pos+process)%64 + 64*((Y-tube_2_Y_Pos)%96)), .data_Out(tube_2_dout));
	  TUBE_3 tube_3_instance(.Clk, .read_address((X-tube_3_X_Pos+process)%64 + 64*((Y-tube_3_Y_Pos)%128)), .data_Out(tube_3_dout));
	  
	  CASTLE castle_instance(.Clk, .read_address((X-castle_X_Pos+process)%160 + 160*((Y-castle_Y_Pos)%160)), .data_Out(castle_dout));
	  
	  STAND stand_instance(.Clk, .read_address((X-Mario_X_Pos+process)%32 + 32*((Y-Mario_Y_Pos)%32)), .data_Out(stand_dout));

//	  BACKGROUND background_instance(.DrawX(X), .DrawY(Y), .process,
//												.cloud_dout, .L_mountain_dout,.S_mountain_dout,.tube_1_dout, .tube_2_dout, .tube_3_dout, .castle_dout,
//												.background_dout,
//												.Cloud_X_Pos, .Cloud_Y_Pos, .L_mountain_X_Pos, .L_mountain_Y_Pos, .S_mountain_X_Pos, .S_mountain_Y_Pos,
//												.tube_1_X_Pos, .tube_1_Y_Pos, .tube_2_X_Pos, .tube_2_Y_Pos, .tube_3_X_Pos, .tube_3_Y_Pos, .castle_X_Pos, .castle_Y_Pos);
	 
	 
	 
	 
	 
	 
	 
	 
    // Display keycode on hex display
    HexDriver hex_inst_0 (keycode[3:0], HEX0);
    HexDriver hex_inst_1 (keycode[7:4], HEX1);
    // HexDriver hex_inst_2 (keycode[11:8], HEX2);
    // HexDriver hex_inst_3 (keycode[15:12], HEX3);
    /**************************************************************************************
        ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
        Hidden Question #1/2:
        What are the advantages and/or disadvantages of using a USB interface over PS/2 interface to
             connect to the keyboard? List any two.  Give an answer in your Post-Lab.
    **************************************************************************************/
endmodule
