//bomb fsm

